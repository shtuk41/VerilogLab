module top_module (
    input clk,
    input a,
    output [3:0] q );
    
    reg [3:0] q_t;
    
    always @(posedge clk) begin
        if (a)
            q_t <= 4'b0100;
        else if (q_t == 4'b0110)
            q_t <= 4'b0000;
        else
            q_t <= q_t + 1'b1;
    end

    assign q = q_t;
    
endmodule
